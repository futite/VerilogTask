`timescale 1ns/1ps
`define DATA_WIDTH  32
`define DATA_DEPTH  1024
`define FIGHT_MODE  3    //可配置为读优先，写优先，保持模式，分别对应为1、2、3
//`define ADDR_WIDTH 10
`define RAM_STYLE_VAL   "block"//"distributed"