`timescale 1ns/1ps
`define  CLK_FREQUENCE  50_000_000
`define  BAUD_RATE       9600
`define  PARITY        "NONE"
`define  FRAME_WD       8
//`define  SAMP_POINT       9