`define DATA_DEPTH 512
`define DATA_WIDTH 32
`define full_min  508
`define empty_max 10
`define FIFO_MODE "Standard"